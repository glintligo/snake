library verilog;
use verilog.vl_types.all;
entity keycheck_vlg_tst is
end keycheck_vlg_tst;

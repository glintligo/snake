library verilog;
use verilog.vl_types.all;
entity random_vlg_tst is
end random_vlg_tst;
